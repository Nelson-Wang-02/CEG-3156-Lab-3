LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY tb_forwardingUnit IS
END tb_forwardingUnit;

ARCHITECTURE testbench OF tb_forwardingUnit IS 

    -- Component Declaration for the Unit Under Test (UUT)
    COMPONENT forwardingUnit
    	port (
			ExMem_RegWrite : IN STD_LOGIC;
			ExMem_Rd, IdEx_Rs, IdEx_Rt : IN STD_LOGIC_VECTOR(4 downto 0);
			
			MemWb_RegWrite : IN STD_LOGIC;
			MemWb_Rd : IN STD_LOGIC_VECTOR(4 downto 0); 
			
			FA1, FA0, FB1, FB0 : OUT STD_LOGIC);
    END COMPONENT;


   --Inputs
   signal tb_EXMEM_RegWrite, tb_MEMWB_RegWrite : STD_LOGIC; 
	signal tb_EXMEM_Rd, tb_IDEX_Rs, tb_IDEX_Rt, tb_MEMWB_Rd : STD_LOGIC_VECTOR(4 downto 0);

    --Outputs
   signal tb_FA1, tb_FA0, tb_FB1, tb_FB0 : STD_LOGIC;

BEGIN 

	-- Instantiate the Unit Under Test (UUT)
   uut: forwardingUnit 
		PORT MAP (
         ExMem_RegWrite => tb_EXMEM_RegWrite,
			ExMem_Rd => tb_EXMEM_Rd, 
			IdEx_Rs => tb_IDEX_Rs, 
			IdEx_Rt => tb_IDEX_Rt,
			
			MemWb_RegWrite => tb_MEMWB_RegWrite,
			MemWb_Rd => tb_MEMWB_Rd,
			
			FA1 => tb_FA1, 
			FA0 => tb_FA0, 
			FB1 => tb_FB1,  
			FB0 => tb_FB0);

   -- Stimulus process
   stim_proc: process
   begin	
      -- hold reset state for 100 ns.
    tb_EXMEM_RegWrite <= '0';
		tb_EXMEM_Rd <= "00000";
		tb_IDEX_Rs <= "00000";
		tb_IDEX_Rt <= "00000";
		tb_MEMWB_RegWrite <= '0';
		tb_MEMWB_Rd <= "00000";
		
		wait for 50 ns;	

		assert tb_FA1 = '0' and tb_FA0 = '0' and tb_FB1 = '0' and tb_FB0 = '0' report "Output should be FA=00 FB=00" severity ERROR; 
		
    tb_EXMEM_RegWrite <= '1';
		tb_EXMEM_Rd <= "00001";
		tb_IDEX_Rs <= "00001";
		tb_IDEX_Rt <= "00001";
		tb_MEMWB_RegWrite <= '0';
		tb_MEMWB_Rd <= "00000";		
		
		wait for 50 ns;	
		
		assert tb_FA1 = '1' and tb_FA0 = '0' and tb_FB1 = '1' and tb_FB0 = '0' report "Output should be FA=10 FB=10" severity ERROR; 
		
    tb_EXMEM_RegWrite <= '0';
		tb_EXMEM_Rd <= "00001";
		tb_IDEX_Rs <= "00001";
		tb_IDEX_Rt <= "00001";
		tb_MEMWB_RegWrite <= '1';
		tb_MEMWB_Rd <= "00001";		
		
		wait for 50 ns;	
		
		assert tb_FA1 = '0' and tb_FA0 = '1' and tb_FB1 = '0' and tb_FB0 = '1' report "Output should be FA=01 FB=01" severity ERROR; 		
      
      wait;
   end process;

END;
